// GitHub thinks the .do files are important and now it thinks the primary language of this repo is "Stata"
// I don't even know what "Stata" is :P

































































































// I hate writing janky things, but I dislike this repo being incorrectly marked as dominantly using "Stata" even more.
