
// change this to change the grid order.
// importing this is not necessary if
// def_griddimensions.sv is imported.
`ifndef DEFINE_GRIDORDER
`define DEFINE_GRIDORDER
    `define GRID_ORD 3
`endif

